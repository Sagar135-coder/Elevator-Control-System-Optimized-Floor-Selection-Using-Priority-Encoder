`timescale 1ns / 1ps
module prioenco_df(d,q);
input [7:0]d;
output [2:0]q;
assign q[2]=~(~(d[7]&d[7])&~(d[6]&d[6])&~(d[5]&d[5])&~(d[4]&d[4]));
assign q[1]=~(~(d[7]&d[7])&~(d[6]&d[6])&~(~(d[5]&d[5])&~(d[4]&d[4])&d[3])&~(~(d[5]&d[5])&~(d[4]&d[4])&d[2]));
assign q[0]=~(~(d[7]&d[7])&~(~(d[6]&d[6])&d[5])&~(~(d[6]&d[6])&~(d[4]&d[4])&d[3])&~(~(d[6]&d[6])&~(d[4]&d[4])&~(d[2]&d[2])&d[1]));
endmodule
